// Controller

module Controller ( opcode,
					funct
					// write your code in here
					);

	input  [5:0] opcode;
    input  [5:0] funct;

	// write your code in here
	
endmodule




